module tb_rom();

//reg clk;
reg [18:0] addr1;
wire [15:0] data1, data2, data3, data4, data5, data6, data7, data8, data9, data10;

rom romp( .addr1(addr1), .data1(data1), .data2(data2), .data3(data3), .data4(data4), .data5(data5),
			 .data6(data6), .data7(data7), .data8(data8), .data9(data9), .data10(data10));


 //always begin
	
  	//clk <=0;
  	//#5;
  	//clk <=1;
	//#5;
  	
  //end

initial begin
//@(negedge clk);
#5 addr1 <= 19'd0;

#5 addr1 <= 19'd10; 

#5 addr1 <= 19'd20;

end
endmodule